library ieee;
use ieee.std_logic_1164.all;

entity test is port(
    data_in, clk : in std_logic;
    data_out : out std_logic;
);
end test;

architecture test_beh of test is

end test_beh;